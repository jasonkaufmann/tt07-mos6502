
module opcode_decoder(
    input [7:0] opcode,
    output reg [3:0] addressing_mode
);

always @(*) begin
    case (opcode)
        8'h00: addressing_mode = 4'b1011;
        8'h01: addressing_mode = 4'b1001;
        8'h05: addressing_mode = 4'b0010;
        8'h06: addressing_mode = 4'b0010;
        8'h08: addressing_mode = 4'b1011;
        8'h09: addressing_mode = 4'b0001;
        8'h0A: addressing_mode = 4'b0000;
        8'h0D: addressing_mode = 4'b0101;
        8'h0E: addressing_mode = 4'b0101;
        8'h10: addressing_mode = 4'b1100;
        8'h11: addressing_mode = 4'b1010;
        8'h15: addressing_mode = 4'b0011;
        8'h16: addressing_mode = 4'b0011;
        8'h18: addressing_mode = 4'b1011;
        8'h19: addressing_mode = 4'b0111;
        8'h1D: addressing_mode = 4'b0110;
        8'h1E: addressing_mode = 4'b0110;
        8'h20: addressing_mode = 4'b0101;
        8'h21: addressing_mode = 4'b1001;
        8'h24: addressing_mode = 4'b0010;
        8'h25: addressing_mode = 4'b0010;
        8'h26: addressing_mode = 4'b0010;
        8'h28: addressing_mode = 4'b1011;
        8'h29: addressing_mode = 4'b0001;
        8'h2A: addressing_mode = 4'b0000;
        8'h2C: addressing_mode = 4'b0101;
        8'h2D: addressing_mode = 4'b0101;
        8'h2E: addressing_mode = 4'b0101;
        8'h30: addressing_mode = 4'b1100;
        8'h31: addressing_mode = 4'b1010;
        8'h35: addressing_mode = 4'b0011;
        8'h36: addressing_mode = 4'b0011;
        8'h38: addressing_mode = 4'b1011;
        8'h39: addressing_mode = 4'b0111;
        8'h3D: addressing_mode = 4'b0110;
        8'h3E: addressing_mode = 4'b0110;
        8'h40: addressing_mode = 4'b1011;
        8'h41: addressing_mode = 4'b1001;
        8'h45: addressing_mode = 4'b0010;
        8'h46: addressing_mode = 4'b0010;
        8'h48: addressing_mode = 4'b1011;
        8'h49: addressing_mode = 4'b0001;
        8'h4A: addressing_mode = 4'b0000;
        8'h4C: addressing_mode = 4'b0101;
        8'h4D: addressing_mode = 4'b0101;
        8'h4E: addressing_mode = 4'b0101;
        8'h50: addressing_mode = 4'b1100;
        8'h51: addressing_mode = 4'b1010;
        8'h55: addressing_mode = 4'b0011;
        8'h56: addressing_mode = 4'b0011;
        8'h58: addressing_mode = 4'b1011;
        8'h59: addressing_mode = 4'b0111;
        8'h5D: addressing_mode = 4'b0110;
        8'h5E: addressing_mode = 4'b0110;
        8'h60: addressing_mode = 4'b1011;
        8'h61: addressing_mode = 4'b1001;
        8'h65: addressing_mode = 4'b0010;
        8'h66: addressing_mode = 4'b0010;
        8'h68: addressing_mode = 4'b1011;
        8'h69: addressing_mode = 4'b0001;
        8'h6A: addressing_mode = 4'b0000;
        8'h6C: addressing_mode = 4'b1000;
        8'h6D: addressing_mode = 4'b0101;
        8'h6E: addressing_mode = 4'b0101;
        8'h70: addressing_mode = 4'b1100;
        8'h71: addressing_mode = 4'b1010;
        8'h75: addressing_mode = 4'b0011;
        8'h76: addressing_mode = 4'b0011;
        8'h78: addressing_mode = 4'b1011;
        8'h79: addressing_mode = 4'b0111;
        8'h7D: addressing_mode = 4'b0110;
        8'h7E: addressing_mode = 4'b0110;
        8'h81: addressing_mode = 4'b1001;
        8'h84: addressing_mode = 4'b0010;
        8'h85: addressing_mode = 4'b0010;
        8'h86: addressing_mode = 4'b0010;
        8'h88: addressing_mode = 4'b1011;
        8'h8A: addressing_mode = 4'b1011;
        8'h8C: addressing_mode = 4'b0101;
        8'h8D: addressing_mode = 4'b0101;
        8'h8E: addressing_mode = 4'b0101;
        8'h90: addressing_mode = 4'b1100;
        8'h91: addressing_mode = 4'b1010;
        8'h94: addressing_mode = 4'b0011;
        8'h95: addressing_mode = 4'b0011;
        8'h96: addressing_mode = 4'b0100;
        8'h98: addressing_mode = 4'b1011;
        8'h99: addressing_mode = 4'b0111;
        8'h9A: addressing_mode = 4'b1011;
        8'h9D: addressing_mode = 4'b0110;
        8'hA0: addressing_mode = 4'b0001;
        8'hA1: addressing_mode = 4'b1001;
        8'hA2: addressing_mode = 4'b0001;
        8'hA4: addressing_mode = 4'b0010;
        8'hA5: addressing_mode = 4'b0010;
        8'hA6: addressing_mode = 4'b0010;
        8'hA8: addressing_mode = 4'b1011;
        8'hA9: addressing_mode = 4'b0001;
        8'hAA: addressing_mode = 4'b1011;
        8'hAC: addressing_mode = 4'b0101;
        8'hAD: addressing_mode = 4'b0101;
        8'hAE: addressing_mode = 4'b0101;
        8'hB0: addressing_mode = 4'b1100;
        8'hB1: addressing_mode = 4'b1010;
        8'hB4: addressing_mode = 4'b0011;
        8'hB5: addressing_mode = 4'b0011;
        8'hB6: addressing_mode = 4'b0100;
        8'hB8: addressing_mode = 4'b1011;
        8'hB9: addressing_mode = 4'b0111;
        8'hBA: addressing_mode = 4'b1011;
        8'hBC: addressing_mode = 4'b0110;
        8'hBD: addressing_mode = 4'b0110;
        8'hBE: addressing_mode = 4'b0111;
        8'hC0: addressing_mode = 4'b0001;
        8'hC1: addressing_mode = 4'b1001;
        8'hC4: addressing_mode = 4'b0010;
        8'hC5: addressing_mode = 4'b0010;
        8'hC6: addressing_mode = 4'b0010;
        8'hC8: addressing_mode = 4'b1011;
        8'hC9: addressing_mode = 4'b0001;
        8'hCA: addressing_mode = 4'b1011;
        8'hCC: addressing_mode = 4'b0101;
        8'hCD: addressing_mode = 4'b0101;
        8'hCE: addressing_mode = 4'b0101;
        8'hD0: addressing_mode = 4'b1100;
        8'hD1: addressing_mode = 4'b1010;
        8'hD5: addressing_mode = 4'b0011;
        8'hD6: addressing_mode = 4'b0011;
        8'hD8: addressing_mode = 4'b1011;
        8'hD9: addressing_mode = 4'b0111;
        8'hDD: addressing_mode = 4'b0110;
        8'hDE: addressing_mode = 4'b0110;
        8'hE0: addressing_mode = 4'b0001;
        8'hE1: addressing_mode = 4'b1001;
        8'hE4: addressing_mode = 4'b0010;
        8'hE5: addressing_mode = 4'b0010;
        8'hE6: addressing_mode = 4'b0010;
        8'hE8: addressing_mode = 4'b1011;
        8'hE9: addressing_mode = 4'b0001;
        8'hEA: addressing_mode = 4'b1011;
        8'hEC: addressing_mode = 4'b0101;
        8'hED: addressing_mode = 4'b0101;
        8'hEE: addressing_mode = 4'b0101;
        8'hF0: addressing_mode = 4'b1100;
        8'hF1: addressing_mode = 4'b1010;
        8'hF5: addressing_mode = 4'b0011;
        8'hF6: addressing_mode = 4'b0011;
        8'hF8: addressing_mode = 4'b1011;
        8'hF9: addressing_mode = 4'b0111;
        8'hFD: addressing_mode = 4'b0110;
        8'hFE: addressing_mode = 4'b0110;

        default: addressing_mode = 4'b1111; // Invalid opcode
    endcase
end

endmodule
